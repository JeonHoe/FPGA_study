library verilog;
use verilog.vl_types.all;
entity tb_de0_memory is
end tb_de0_memory;
