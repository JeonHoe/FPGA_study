library verilog;
use verilog.vl_types.all;
entity tb_final is
end tb_final;
