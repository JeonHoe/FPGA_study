library verilog;
use verilog.vl_types.all;
entity tb_de0_doorlock_fixed is
end tb_de0_doorlock_fixed;
